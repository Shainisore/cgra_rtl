typedef struct packed {
  logic [5:0] ctrl ;
  logic [0:0] predicate ;
  logic [3:0][2:0] fu_in ;
  logic [7:0][2:0] outport ;
  logic [5:0][0:0] predicate_in ;
} CGRAConfig_6_4_6_8;

typedef struct packed {
  logic [31:0] payload ;
  logic [0:0] predicate ;
  logic [0:0] bypass ;
} CGRAData_32_1_1;

typedef struct packed {
  logic [0:0] payload ;
  logic [0:0] predicate ;
} CGRAData_1_1;

module top
(
  input logic [0:0] clk,
  input logic [0:0] reset,
  input logic [0:0] recv_waddr__en [0:15],
  input logic [1:0] recv_waddr__msg [0:15],
  output logic [0:0] recv_waddr__rdy [0:15],
  input logic [0:0] recv_wopt__en [0:15],
  input CGRAConfig_6_4_6_8 recv_wopt__msg [0:15],
  output logic [0:0] recv_wopt__rdy [0:15]
);
  //-------------------------------------------------------------
  // Component data_mem
  //-------------------------------------------------------------

  logic [0:0] data_mem__clk ;
  logic [0:0] data_mem__reset ;
  logic [0:0] data_mem__recv_raddr__en [0:3] ;
  logic [6:0] data_mem__recv_raddr__msg [0:3] ;
  logic [0:0] data_mem__recv_raddr__rdy [0:3] ;
  logic [0:0] data_mem__recv_waddr__en [0:3] ;
  logic [6:0] data_mem__recv_waddr__msg [0:3] ;
  logic [0:0] data_mem__recv_waddr__rdy [0:3] ;
  logic [0:0] data_mem__recv_wdata__en [0:3] ;
  CGRAData_32_1_1 data_mem__recv_wdata__msg [0:3] ;
  logic [0:0] data_mem__recv_wdata__rdy [0:3] ;
  logic [0:0] data_mem__send_rdata__en [0:3] ;
  CGRAData_32_1_1 data_mem__send_rdata__msg [0:3] ;
  logic [0:0] data_mem__send_rdata__rdy [0:3] ;

  DataMemRTL__2aacae905ddf1f6e data_mem
  (
    .clk( data_mem__clk ),
    .reset( data_mem__reset ),
    .recv_raddr__en( data_mem__recv_raddr__en ),
    .recv_raddr__msg( data_mem__recv_raddr__msg ),
    .recv_raddr__rdy( data_mem__recv_raddr__rdy ),
    .recv_waddr__en( data_mem__recv_waddr__en ),
    .recv_waddr__msg( data_mem__recv_waddr__msg ),
    .recv_waddr__rdy( data_mem__recv_waddr__rdy ),
    .recv_wdata__en( data_mem__recv_wdata__en ),
    .recv_wdata__msg( data_mem__recv_wdata__msg ),
    .recv_wdata__rdy( data_mem__recv_wdata__rdy ),
    .send_rdata__en( data_mem__send_rdata__en ),
    .send_rdata__msg( data_mem__send_rdata__msg ),
    .send_rdata__rdy( data_mem__send_rdata__rdy )
  );

  //-------------------------------------------------------------
  // End of component data_mem
  //-------------------------------------------------------------

  //-------------------------------------------------------------
  // Component tile[0:15]
  //-------------------------------------------------------------

  logic [0:0] tile__clk [0:15] ;
  logic [0:0] tile__reset [0:15] ;
  logic [0:0] tile__from_mem_rdata__en [0:15] ;
  CGRAData_32_1_1 tile__from_mem_rdata__msg [0:15] ;
  logic [0:0] tile__from_mem_rdata__rdy [0:15] ;
  logic [0:0] tile__recv_data__en [0:15][0:3] ;
  CGRAData_32_1_1 tile__recv_data__msg [0:15][0:3] ;
  logic [0:0] tile__recv_data__rdy [0:15][0:3] ;
  logic [0:0] tile__recv_waddr__en [0:15] ;
  logic [1:0] tile__recv_waddr__msg [0:15] ;
  logic [0:0] tile__recv_waddr__rdy [0:15] ;
  logic [0:0] tile__recv_wopt__en [0:15] ;
  CGRAConfig_6_4_6_8 tile__recv_wopt__msg [0:15] ;
  logic [0:0] tile__recv_wopt__rdy [0:15] ;
  logic [0:0] tile__send_data__en [0:15][0:3] ;
  CGRAData_32_1_1 tile__send_data__msg [0:15][0:3] ;
  logic [0:0] tile__send_data__rdy [0:15][0:3] ;
  logic [0:0] tile__to_mem_raddr__en [0:15] ;
  logic [6:0] tile__to_mem_raddr__msg [0:15] ;
  logic [0:0] tile__to_mem_raddr__rdy [0:15] ;
  logic [0:0] tile__to_mem_waddr__en [0:15] ;
  logic [6:0] tile__to_mem_waddr__msg [0:15] ;
  logic [0:0] tile__to_mem_waddr__rdy [0:15] ;
  logic [0:0] tile__to_mem_wdata__en [0:15] ;
  CGRAData_32_1_1 tile__to_mem_wdata__msg [0:15] ;
  logic [0:0] tile__to_mem_wdata__rdy [0:15] ;

  TileRTL__97e625cd3d6bdc66 tile__0
  (
    .clk( tile__clk[0] ),
    .reset( tile__reset[0] ),
    .from_mem_rdata__en( tile__from_mem_rdata__en[0] ),
    .from_mem_rdata__msg( tile__from_mem_rdata__msg[0] ),
    .from_mem_rdata__rdy( tile__from_mem_rdata__rdy[0] ),
    .recv_data__en( tile__recv_data__en[0] ),
    .recv_data__msg( tile__recv_data__msg[0] ),
    .recv_data__rdy( tile__recv_data__rdy[0] ),
    .recv_waddr__en( tile__recv_waddr__en[0] ),
    .recv_waddr__msg( tile__recv_waddr__msg[0] ),
    .recv_waddr__rdy( tile__recv_waddr__rdy[0] ),
    .recv_wopt__en( tile__recv_wopt__en[0] ),
    .recv_wopt__msg( tile__recv_wopt__msg[0] ),
    .recv_wopt__rdy( tile__recv_wopt__rdy[0] ),
    .send_data__en( tile__send_data__en[0] ),
    .send_data__msg( tile__send_data__msg[0] ),
    .send_data__rdy( tile__send_data__rdy[0] ),
    .to_mem_raddr__en( tile__to_mem_raddr__en[0] ),
    .to_mem_raddr__msg( tile__to_mem_raddr__msg[0] ),
    .to_mem_raddr__rdy( tile__to_mem_raddr__rdy[0] ),
    .to_mem_waddr__en( tile__to_mem_waddr__en[0] ),
    .to_mem_waddr__msg( tile__to_mem_waddr__msg[0] ),
    .to_mem_waddr__rdy( tile__to_mem_waddr__rdy[0] ),
    .to_mem_wdata__en( tile__to_mem_wdata__en[0] ),
    .to_mem_wdata__msg( tile__to_mem_wdata__msg[0] ),
    .to_mem_wdata__rdy( tile__to_mem_wdata__rdy[0] )
  );

  TileRTL__97e625cd3d6bdc66 tile__1
  (
    .clk( tile__clk[1] ),
    .reset( tile__reset[1] ),
    .from_mem_rdata__en( tile__from_mem_rdata__en[1] ),
    .from_mem_rdata__msg( tile__from_mem_rdata__msg[1] ),
    .from_mem_rdata__rdy( tile__from_mem_rdata__rdy[1] ),
    .recv_data__en( tile__recv_data__en[1] ),
    .recv_data__msg( tile__recv_data__msg[1] ),
    .recv_data__rdy( tile__recv_data__rdy[1] ),
    .recv_waddr__en( tile__recv_waddr__en[1] ),
    .recv_waddr__msg( tile__recv_waddr__msg[1] ),
    .recv_waddr__rdy( tile__recv_waddr__rdy[1] ),
    .recv_wopt__en( tile__recv_wopt__en[1] ),
    .recv_wopt__msg( tile__recv_wopt__msg[1] ),
    .recv_wopt__rdy( tile__recv_wopt__rdy[1] ),
    .send_data__en( tile__send_data__en[1] ),
    .send_data__msg( tile__send_data__msg[1] ),
    .send_data__rdy( tile__send_data__rdy[1] ),
    .to_mem_raddr__en( tile__to_mem_raddr__en[1] ),
    .to_mem_raddr__msg( tile__to_mem_raddr__msg[1] ),
    .to_mem_raddr__rdy( tile__to_mem_raddr__rdy[1] ),
    .to_mem_waddr__en( tile__to_mem_waddr__en[1] ),
    .to_mem_waddr__msg( tile__to_mem_waddr__msg[1] ),
    .to_mem_waddr__rdy( tile__to_mem_waddr__rdy[1] ),
    .to_mem_wdata__en( tile__to_mem_wdata__en[1] ),
    .to_mem_wdata__msg( tile__to_mem_wdata__msg[1] ),
    .to_mem_wdata__rdy( tile__to_mem_wdata__rdy[1] )
  );

  TileRTL__97e625cd3d6bdc66 tile__2
  (
    .clk( tile__clk[2] ),
    .reset( tile__reset[2] ),
    .from_mem_rdata__en( tile__from_mem_rdata__en[2] ),
    .from_mem_rdata__msg( tile__from_mem_rdata__msg[2] ),
    .from_mem_rdata__rdy( tile__from_mem_rdata__rdy[2] ),
    .recv_data__en( tile__recv_data__en[2] ),
    .recv_data__msg( tile__recv_data__msg[2] ),
    .recv_data__rdy( tile__recv_data__rdy[2] ),
    .recv_waddr__en( tile__recv_waddr__en[2] ),
    .recv_waddr__msg( tile__recv_waddr__msg[2] ),
    .recv_waddr__rdy( tile__recv_waddr__rdy[2] ),
    .recv_wopt__en( tile__recv_wopt__en[2] ),
    .recv_wopt__msg( tile__recv_wopt__msg[2] ),
    .recv_wopt__rdy( tile__recv_wopt__rdy[2] ),
    .send_data__en( tile__send_data__en[2] ),
    .send_data__msg( tile__send_data__msg[2] ),
    .send_data__rdy( tile__send_data__rdy[2] ),
    .to_mem_raddr__en( tile__to_mem_raddr__en[2] ),
    .to_mem_raddr__msg( tile__to_mem_raddr__msg[2] ),
    .to_mem_raddr__rdy( tile__to_mem_raddr__rdy[2] ),
    .to_mem_waddr__en( tile__to_mem_waddr__en[2] ),
    .to_mem_waddr__msg( tile__to_mem_waddr__msg[2] ),
    .to_mem_waddr__rdy( tile__to_mem_waddr__rdy[2] ),
    .to_mem_wdata__en( tile__to_mem_wdata__en[2] ),
    .to_mem_wdata__msg( tile__to_mem_wdata__msg[2] ),
    .to_mem_wdata__rdy( tile__to_mem_wdata__rdy[2] )
  );

  TileRTL__97e625cd3d6bdc66 tile__3
  (
    .clk( tile__clk[3] ),
    .reset( tile__reset[3] ),
    .from_mem_rdata__en( tile__from_mem_rdata__en[3] ),
    .from_mem_rdata__msg( tile__from_mem_rdata__msg[3] ),
    .from_mem_rdata__rdy( tile__from_mem_rdata__rdy[3] ),
    .recv_data__en( tile__recv_data__en[3] ),
    .recv_data__msg( tile__recv_data__msg[3] ),
    .recv_data__rdy( tile__recv_data__rdy[3] ),
    .recv_waddr__en( tile__recv_waddr__en[3] ),
    .recv_waddr__msg( tile__recv_waddr__msg[3] ),
    .recv_waddr__rdy( tile__recv_waddr__rdy[3] ),
    .recv_wopt__en( tile__recv_wopt__en[3] ),
    .recv_wopt__msg( tile__recv_wopt__msg[3] ),
    .recv_wopt__rdy( tile__recv_wopt__rdy[3] ),
    .send_data__en( tile__send_data__en[3] ),
    .send_data__msg( tile__send_data__msg[3] ),
    .send_data__rdy( tile__send_data__rdy[3] ),
    .to_mem_raddr__en( tile__to_mem_raddr__en[3] ),
    .to_mem_raddr__msg( tile__to_mem_raddr__msg[3] ),
    .to_mem_raddr__rdy( tile__to_mem_raddr__rdy[3] ),
    .to_mem_waddr__en( tile__to_mem_waddr__en[3] ),
    .to_mem_waddr__msg( tile__to_mem_waddr__msg[3] ),
    .to_mem_waddr__rdy( tile__to_mem_waddr__rdy[3] ),
    .to_mem_wdata__en( tile__to_mem_wdata__en[3] ),
    .to_mem_wdata__msg( tile__to_mem_wdata__msg[3] ),
    .to_mem_wdata__rdy( tile__to_mem_wdata__rdy[3] )
  );

  TileRTL__97e625cd3d6bdc66 tile__4
  (
    .clk( tile__clk[4] ),
    .reset( tile__reset[4] ),
    .from_mem_rdata__en( tile__from_mem_rdata__en[4] ),
    .from_mem_rdata__msg( tile__from_mem_rdata__msg[4] ),
    .from_mem_rdata__rdy( tile__from_mem_rdata__rdy[4] ),
    .recv_data__en( tile__recv_data__en[4] ),
    .recv_data__msg( tile__recv_data__msg[4] ),
    .recv_data__rdy( tile__recv_data__rdy[4] ),
    .recv_waddr__en( tile__recv_waddr__en[4] ),
    .recv_waddr__msg( tile__recv_waddr__msg[4] ),
    .recv_waddr__rdy( tile__recv_waddr__rdy[4] ),
    .recv_wopt__en( tile__recv_wopt__en[4] ),
    .recv_wopt__msg( tile__recv_wopt__msg[4] ),
    .recv_wopt__rdy( tile__recv_wopt__rdy[4] ),
    .send_data__en( tile__send_data__en[4] ),
    .send_data__msg( tile__send_data__msg[4] ),
    .send_data__rdy( tile__send_data__rdy[4] ),
    .to_mem_raddr__en( tile__to_mem_raddr__en[4] ),
    .to_mem_raddr__msg( tile__to_mem_raddr__msg[4] ),
    .to_mem_raddr__rdy( tile__to_mem_raddr__rdy[4] ),
    .to_mem_waddr__en( tile__to_mem_waddr__en[4] ),
    .to_mem_waddr__msg( tile__to_mem_waddr__msg[4] ),
    .to_mem_waddr__rdy( tile__to_mem_waddr__rdy[4] ),
    .to_mem_wdata__en( tile__to_mem_wdata__en[4] ),
    .to_mem_wdata__msg( tile__to_mem_wdata__msg[4] ),
    .to_mem_wdata__rdy( tile__to_mem_wdata__rdy[4] )
  );

  TileRTL__97e625cd3d6bdc66 tile__5
  (
    .clk( tile__clk[5] ),
    .reset( tile__reset[5] ),
    .from_mem_rdata__en( tile__from_mem_rdata__en[5] ),
    .from_mem_rdata__msg( tile__from_mem_rdata__msg[5] ),
    .from_mem_rdata__rdy( tile__from_mem_rdata__rdy[5] ),
    .recv_data__en( tile__recv_data__en[5] ),
    .recv_data__msg( tile__recv_data__msg[5] ),
    .recv_data__rdy( tile__recv_data__rdy[5] ),
    .recv_waddr__en( tile__recv_waddr__en[5] ),
    .recv_waddr__msg( tile__recv_waddr__msg[5] ),
    .recv_waddr__rdy( tile__recv_waddr__rdy[5] ),
    .recv_wopt__en( tile__recv_wopt__en[5] ),
    .recv_wopt__msg( tile__recv_wopt__msg[5] ),
    .recv_wopt__rdy( tile__recv_wopt__rdy[5] ),
    .send_data__en( tile__send_data__en[5] ),
    .send_data__msg( tile__send_data__msg[5] ),
    .send_data__rdy( tile__send_data__rdy[5] ),
    .to_mem_raddr__en( tile__to_mem_raddr__en[5] ),
    .to_mem_raddr__msg( tile__to_mem_raddr__msg[5] ),
    .to_mem_raddr__rdy( tile__to_mem_raddr__rdy[5] ),
    .to_mem_waddr__en( tile__to_mem_waddr__en[5] ),
    .to_mem_waddr__msg( tile__to_mem_waddr__msg[5] ),
    .to_mem_waddr__rdy( tile__to_mem_waddr__rdy[5] ),
    .to_mem_wdata__en( tile__to_mem_wdata__en[5] ),
    .to_mem_wdata__msg( tile__to_mem_wdata__msg[5] ),
    .to_mem_wdata__rdy( tile__to_mem_wdata__rdy[5] )
  );

  TileRTL__97e625cd3d6bdc66 tile__6
  (
    .clk( tile__clk[6] ),
    .reset( tile__reset[6] ),
    .from_mem_rdata__en( tile__from_mem_rdata__en[6] ),
    .from_mem_rdata__msg( tile__from_mem_rdata__msg[6] ),
    .from_mem_rdata__rdy( tile__from_mem_rdata__rdy[6] ),
    .recv_data__en( tile__recv_data__en[6] ),
    .recv_data__msg( tile__recv_data__msg[6] ),
    .recv_data__rdy( tile__recv_data__rdy[6] ),
    .recv_waddr__en( tile__recv_waddr__en[6] ),
    .recv_waddr__msg( tile__recv_waddr__msg[6] ),
    .recv_waddr__rdy( tile__recv_waddr__rdy[6] ),
    .recv_wopt__en( tile__recv_wopt__en[6] ),
    .recv_wopt__msg( tile__recv_wopt__msg[6] ),
    .recv_wopt__rdy( tile__recv_wopt__rdy[6] ),
    .send_data__en( tile__send_data__en[6] ),
    .send_data__msg( tile__send_data__msg[6] ),
    .send_data__rdy( tile__send_data__rdy[6] ),
    .to_mem_raddr__en( tile__to_mem_raddr__en[6] ),
    .to_mem_raddr__msg( tile__to_mem_raddr__msg[6] ),
    .to_mem_raddr__rdy( tile__to_mem_raddr__rdy[6] ),
    .to_mem_waddr__en( tile__to_mem_waddr__en[6] ),
    .to_mem_waddr__msg( tile__to_mem_waddr__msg[6] ),
    .to_mem_waddr__rdy( tile__to_mem_waddr__rdy[6] ),
    .to_mem_wdata__en( tile__to_mem_wdata__en[6] ),
    .to_mem_wdata__msg( tile__to_mem_wdata__msg[6] ),
    .to_mem_wdata__rdy( tile__to_mem_wdata__rdy[6] )
  );

  TileRTL__97e625cd3d6bdc66 tile__7
  (
    .clk( tile__clk[7] ),
    .reset( tile__reset[7] ),
    .from_mem_rdata__en( tile__from_mem_rdata__en[7] ),
    .from_mem_rdata__msg( tile__from_mem_rdata__msg[7] ),
    .from_mem_rdata__rdy( tile__from_mem_rdata__rdy[7] ),
    .recv_data__en( tile__recv_data__en[7] ),
    .recv_data__msg( tile__recv_data__msg[7] ),
    .recv_data__rdy( tile__recv_data__rdy[7] ),
    .recv_waddr__en( tile__recv_waddr__en[7] ),
    .recv_waddr__msg( tile__recv_waddr__msg[7] ),
    .recv_waddr__rdy( tile__recv_waddr__rdy[7] ),
    .recv_wopt__en( tile__recv_wopt__en[7] ),
    .recv_wopt__msg( tile__recv_wopt__msg[7] ),
    .recv_wopt__rdy( tile__recv_wopt__rdy[7] ),
    .send_data__en( tile__send_data__en[7] ),
    .send_data__msg( tile__send_data__msg[7] ),
    .send_data__rdy( tile__send_data__rdy[7] ),
    .to_mem_raddr__en( tile__to_mem_raddr__en[7] ),
    .to_mem_raddr__msg( tile__to_mem_raddr__msg[7] ),
    .to_mem_raddr__rdy( tile__to_mem_raddr__rdy[7] ),
    .to_mem_waddr__en( tile__to_mem_waddr__en[7] ),
    .to_mem_waddr__msg( tile__to_mem_waddr__msg[7] ),
    .to_mem_waddr__rdy( tile__to_mem_waddr__rdy[7] ),
    .to_mem_wdata__en( tile__to_mem_wdata__en[7] ),
    .to_mem_wdata__msg( tile__to_mem_wdata__msg[7] ),
    .to_mem_wdata__rdy( tile__to_mem_wdata__rdy[7] )
  );

  TileRTL__97e625cd3d6bdc66 tile__8
  (
    .clk( tile__clk[8] ),
    .reset( tile__reset[8] ),
    .from_mem_rdata__en( tile__from_mem_rdata__en[8] ),
    .from_mem_rdata__msg( tile__from_mem_rdata__msg[8] ),
    .from_mem_rdata__rdy( tile__from_mem_rdata__rdy[8] ),
    .recv_data__en( tile__recv_data__en[8] ),
    .recv_data__msg( tile__recv_data__msg[8] ),
    .recv_data__rdy( tile__recv_data__rdy[8] ),
    .recv_waddr__en( tile__recv_waddr__en[8] ),
    .recv_waddr__msg( tile__recv_waddr__msg[8] ),
    .recv_waddr__rdy( tile__recv_waddr__rdy[8] ),
    .recv_wopt__en( tile__recv_wopt__en[8] ),
    .recv_wopt__msg( tile__recv_wopt__msg[8] ),
    .recv_wopt__rdy( tile__recv_wopt__rdy[8] ),
    .send_data__en( tile__send_data__en[8] ),
    .send_data__msg( tile__send_data__msg[8] ),
    .send_data__rdy( tile__send_data__rdy[8] ),
    .to_mem_raddr__en( tile__to_mem_raddr__en[8] ),
    .to_mem_raddr__msg( tile__to_mem_raddr__msg[8] ),
    .to_mem_raddr__rdy( tile__to_mem_raddr__rdy[8] ),
    .to_mem_waddr__en( tile__to_mem_waddr__en[8] ),
    .to_mem_waddr__msg( tile__to_mem_waddr__msg[8] ),
    .to_mem_waddr__rdy( tile__to_mem_waddr__rdy[8] ),
    .to_mem_wdata__en( tile__to_mem_wdata__en[8] ),
    .to_mem_wdata__msg( tile__to_mem_wdata__msg[8] ),
    .to_mem_wdata__rdy( tile__to_mem_wdata__rdy[8] )
  );

  TileRTL__97e625cd3d6bdc66 tile__9
  (
    .clk( tile__clk[9] ),
    .reset( tile__reset[9] ),
    .from_mem_rdata__en( tile__from_mem_rdata__en[9] ),
    .from_mem_rdata__msg( tile__from_mem_rdata__msg[9] ),
    .from_mem_rdata__rdy( tile__from_mem_rdata__rdy[9] ),
    .recv_data__en( tile__recv_data__en[9] ),
    .recv_data__msg( tile__recv_data__msg[9] ),
    .recv_data__rdy( tile__recv_data__rdy[9] ),
    .recv_waddr__en( tile__recv_waddr__en[9] ),
    .recv_waddr__msg( tile__recv_waddr__msg[9] ),
    .recv_waddr__rdy( tile__recv_waddr__rdy[9] ),
    .recv_wopt__en( tile__recv_wopt__en[9] ),
    .recv_wopt__msg( tile__recv_wopt__msg[9] ),
    .recv_wopt__rdy( tile__recv_wopt__rdy[9] ),
    .send_data__en( tile__send_data__en[9] ),
    .send_data__msg( tile__send_data__msg[9] ),
    .send_data__rdy( tile__send_data__rdy[9] ),
    .to_mem_raddr__en( tile__to_mem_raddr__en[9] ),
    .to_mem_raddr__msg( tile__to_mem_raddr__msg[9] ),
    .to_mem_raddr__rdy( tile__to_mem_raddr__rdy[9] ),
    .to_mem_waddr__en( tile__to_mem_waddr__en[9] ),
    .to_mem_waddr__msg( tile__to_mem_waddr__msg[9] ),
    .to_mem_waddr__rdy( tile__to_mem_waddr__rdy[9] ),
    .to_mem_wdata__en( tile__to_mem_wdata__en[9] ),
    .to_mem_wdata__msg( tile__to_mem_wdata__msg[9] ),
    .to_mem_wdata__rdy( tile__to_mem_wdata__rdy[9] )
  );

  TileRTL__97e625cd3d6bdc66 tile__10
  (
    .clk( tile__clk[10] ),
    .reset( tile__reset[10] ),
    .from_mem_rdata__en( tile__from_mem_rdata__en[10] ),
    .from_mem_rdata__msg( tile__from_mem_rdata__msg[10] ),
    .from_mem_rdata__rdy( tile__from_mem_rdata__rdy[10] ),
    .recv_data__en( tile__recv_data__en[10] ),
    .recv_data__msg( tile__recv_data__msg[10] ),
    .recv_data__rdy( tile__recv_data__rdy[10] ),
    .recv_waddr__en( tile__recv_waddr__en[10] ),
    .recv_waddr__msg( tile__recv_waddr__msg[10] ),
    .recv_waddr__rdy( tile__recv_waddr__rdy[10] ),
    .recv_wopt__en( tile__recv_wopt__en[10] ),
    .recv_wopt__msg( tile__recv_wopt__msg[10] ),
    .recv_wopt__rdy( tile__recv_wopt__rdy[10] ),
    .send_data__en( tile__send_data__en[10] ),
    .send_data__msg( tile__send_data__msg[10] ),
    .send_data__rdy( tile__send_data__rdy[10] ),
    .to_mem_raddr__en( tile__to_mem_raddr__en[10] ),
    .to_mem_raddr__msg( tile__to_mem_raddr__msg[10] ),
    .to_mem_raddr__rdy( tile__to_mem_raddr__rdy[10] ),
    .to_mem_waddr__en( tile__to_mem_waddr__en[10] ),
    .to_mem_waddr__msg( tile__to_mem_waddr__msg[10] ),
    .to_mem_waddr__rdy( tile__to_mem_waddr__rdy[10] ),
    .to_mem_wdata__en( tile__to_mem_wdata__en[10] ),
    .to_mem_wdata__msg( tile__to_mem_wdata__msg[10] ),
    .to_mem_wdata__rdy( tile__to_mem_wdata__rdy[10] )
  );

  TileRTL__97e625cd3d6bdc66 tile__11
  (
    .clk( tile__clk[11] ),
    .reset( tile__reset[11] ),
    .from_mem_rdata__en( tile__from_mem_rdata__en[11] ),
    .from_mem_rdata__msg( tile__from_mem_rdata__msg[11] ),
    .from_mem_rdata__rdy( tile__from_mem_rdata__rdy[11] ),
    .recv_data__en( tile__recv_data__en[11] ),
    .recv_data__msg( tile__recv_data__msg[11] ),
    .recv_data__rdy( tile__recv_data__rdy[11] ),
    .recv_waddr__en( tile__recv_waddr__en[11] ),
    .recv_waddr__msg( tile__recv_waddr__msg[11] ),
    .recv_waddr__rdy( tile__recv_waddr__rdy[11] ),
    .recv_wopt__en( tile__recv_wopt__en[11] ),
    .recv_wopt__msg( tile__recv_wopt__msg[11] ),
    .recv_wopt__rdy( tile__recv_wopt__rdy[11] ),
    .send_data__en( tile__send_data__en[11] ),
    .send_data__msg( tile__send_data__msg[11] ),
    .send_data__rdy( tile__send_data__rdy[11] ),
    .to_mem_raddr__en( tile__to_mem_raddr__en[11] ),
    .to_mem_raddr__msg( tile__to_mem_raddr__msg[11] ),
    .to_mem_raddr__rdy( tile__to_mem_raddr__rdy[11] ),
    .to_mem_waddr__en( tile__to_mem_waddr__en[11] ),
    .to_mem_waddr__msg( tile__to_mem_waddr__msg[11] ),
    .to_mem_waddr__rdy( tile__to_mem_waddr__rdy[11] ),
    .to_mem_wdata__en( tile__to_mem_wdata__en[11] ),
    .to_mem_wdata__msg( tile__to_mem_wdata__msg[11] ),
    .to_mem_wdata__rdy( tile__to_mem_wdata__rdy[11] )
  );

  TileRTL__97e625cd3d6bdc66 tile__12
  (
    .clk( tile__clk[12] ),
    .reset( tile__reset[12] ),
    .from_mem_rdata__en( tile__from_mem_rdata__en[12] ),
    .from_mem_rdata__msg( tile__from_mem_rdata__msg[12] ),
    .from_mem_rdata__rdy( tile__from_mem_rdata__rdy[12] ),
    .recv_data__en( tile__recv_data__en[12] ),
    .recv_data__msg( tile__recv_data__msg[12] ),
    .recv_data__rdy( tile__recv_data__rdy[12] ),
    .recv_waddr__en( tile__recv_waddr__en[12] ),
    .recv_waddr__msg( tile__recv_waddr__msg[12] ),
    .recv_waddr__rdy( tile__recv_waddr__rdy[12] ),
    .recv_wopt__en( tile__recv_wopt__en[12] ),
    .recv_wopt__msg( tile__recv_wopt__msg[12] ),
    .recv_wopt__rdy( tile__recv_wopt__rdy[12] ),
    .send_data__en( tile__send_data__en[12] ),
    .send_data__msg( tile__send_data__msg[12] ),
    .send_data__rdy( tile__send_data__rdy[12] ),
    .to_mem_raddr__en( tile__to_mem_raddr__en[12] ),
    .to_mem_raddr__msg( tile__to_mem_raddr__msg[12] ),
    .to_mem_raddr__rdy( tile__to_mem_raddr__rdy[12] ),
    .to_mem_waddr__en( tile__to_mem_waddr__en[12] ),
    .to_mem_waddr__msg( tile__to_mem_waddr__msg[12] ),
    .to_mem_waddr__rdy( tile__to_mem_waddr__rdy[12] ),
    .to_mem_wdata__en( tile__to_mem_wdata__en[12] ),
    .to_mem_wdata__msg( tile__to_mem_wdata__msg[12] ),
    .to_mem_wdata__rdy( tile__to_mem_wdata__rdy[12] )
  );

  TileRTL__97e625cd3d6bdc66 tile__13
  (
    .clk( tile__clk[13] ),
    .reset( tile__reset[13] ),
    .from_mem_rdata__en( tile__from_mem_rdata__en[13] ),
    .from_mem_rdata__msg( tile__from_mem_rdata__msg[13] ),
    .from_mem_rdata__rdy( tile__from_mem_rdata__rdy[13] ),
    .recv_data__en( tile__recv_data__en[13] ),
    .recv_data__msg( tile__recv_data__msg[13] ),
    .recv_data__rdy( tile__recv_data__rdy[13] ),
    .recv_waddr__en( tile__recv_waddr__en[13] ),
    .recv_waddr__msg( tile__recv_waddr__msg[13] ),
    .recv_waddr__rdy( tile__recv_waddr__rdy[13] ),
    .recv_wopt__en( tile__recv_wopt__en[13] ),
    .recv_wopt__msg( tile__recv_wopt__msg[13] ),
    .recv_wopt__rdy( tile__recv_wopt__rdy[13] ),
    .send_data__en( tile__send_data__en[13] ),
    .send_data__msg( tile__send_data__msg[13] ),
    .send_data__rdy( tile__send_data__rdy[13] ),
    .to_mem_raddr__en( tile__to_mem_raddr__en[13] ),
    .to_mem_raddr__msg( tile__to_mem_raddr__msg[13] ),
    .to_mem_raddr__rdy( tile__to_mem_raddr__rdy[13] ),
    .to_mem_waddr__en( tile__to_mem_waddr__en[13] ),
    .to_mem_waddr__msg( tile__to_mem_waddr__msg[13] ),
    .to_mem_waddr__rdy( tile__to_mem_waddr__rdy[13] ),
    .to_mem_wdata__en( tile__to_mem_wdata__en[13] ),
    .to_mem_wdata__msg( tile__to_mem_wdata__msg[13] ),
    .to_mem_wdata__rdy( tile__to_mem_wdata__rdy[13] )
  );

  TileRTL__97e625cd3d6bdc66 tile__14
  (
    .clk( tile__clk[14] ),
    .reset( tile__reset[14] ),
    .from_mem_rdata__en( tile__from_mem_rdata__en[14] ),
    .from_mem_rdata__msg( tile__from_mem_rdata__msg[14] ),
    .from_mem_rdata__rdy( tile__from_mem_rdata__rdy[14] ),
    .recv_data__en( tile__recv_data__en[14] ),
    .recv_data__msg( tile__recv_data__msg[14] ),
    .recv_data__rdy( tile__recv_data__rdy[14] ),
    .recv_waddr__en( tile__recv_waddr__en[14] ),
    .recv_waddr__msg( tile__recv_waddr__msg[14] ),
    .recv_waddr__rdy( tile__recv_waddr__rdy[14] ),
    .recv_wopt__en( tile__recv_wopt__en[14] ),
    .recv_wopt__msg( tile__recv_wopt__msg[14] ),
    .recv_wopt__rdy( tile__recv_wopt__rdy[14] ),
    .send_data__en( tile__send_data__en[14] ),
    .send_data__msg( tile__send_data__msg[14] ),
    .send_data__rdy( tile__send_data__rdy[14] ),
    .to_mem_raddr__en( tile__to_mem_raddr__en[14] ),
    .to_mem_raddr__msg( tile__to_mem_raddr__msg[14] ),
    .to_mem_raddr__rdy( tile__to_mem_raddr__rdy[14] ),
    .to_mem_waddr__en( tile__to_mem_waddr__en[14] ),
    .to_mem_waddr__msg( tile__to_mem_waddr__msg[14] ),
    .to_mem_waddr__rdy( tile__to_mem_waddr__rdy[14] ),
    .to_mem_wdata__en( tile__to_mem_wdata__en[14] ),
    .to_mem_wdata__msg( tile__to_mem_wdata__msg[14] ),
    .to_mem_wdata__rdy( tile__to_mem_wdata__rdy[14] )
  );

  TileRTL__97e625cd3d6bdc66 tile__15
  (
    .clk( tile__clk[15] ),
    .reset( tile__reset[15] ),
    .from_mem_rdata__en( tile__from_mem_rdata__en[15] ),
    .from_mem_rdata__msg( tile__from_mem_rdata__msg[15] ),
    .from_mem_rdata__rdy( tile__from_mem_rdata__rdy[15] ),
    .recv_data__en( tile__recv_data__en[15] ),
    .recv_data__msg( tile__recv_data__msg[15] ),
    .recv_data__rdy( tile__recv_data__rdy[15] ),
    .recv_waddr__en( tile__recv_waddr__en[15] ),
    .recv_waddr__msg( tile__recv_waddr__msg[15] ),
    .recv_waddr__rdy( tile__recv_waddr__rdy[15] ),
    .recv_wopt__en( tile__recv_wopt__en[15] ),
    .recv_wopt__msg( tile__recv_wopt__msg[15] ),
    .recv_wopt__rdy( tile__recv_wopt__rdy[15] ),
    .send_data__en( tile__send_data__en[15] ),
    .send_data__msg( tile__send_data__msg[15] ),
    .send_data__rdy( tile__send_data__rdy[15] ),
    .to_mem_raddr__en( tile__to_mem_raddr__en[15] ),
    .to_mem_raddr__msg( tile__to_mem_raddr__msg[15] ),
    .to_mem_raddr__rdy( tile__to_mem_raddr__rdy[15] ),
    .to_mem_waddr__en( tile__to_mem_waddr__en[15] ),
    .to_mem_waddr__msg( tile__to_mem_waddr__msg[15] ),
    .to_mem_waddr__rdy( tile__to_mem_waddr__rdy[15] ),
    .to_mem_wdata__en( tile__to_mem_wdata__en[15] ),
    .to_mem_wdata__msg( tile__to_mem_wdata__msg[15] ),
    .to_mem_wdata__rdy( tile__to_mem_wdata__rdy[15] )
  );

  //-------------------------------------------------------------
  // End of component tile[0:15]
  //-------------------------------------------------------------

  assign tile__clk[0] = clk;
  assign tile__reset[0] = reset;
  assign tile__clk[1] = clk;
  assign tile__reset[1] = reset;
  assign tile__clk[2] = clk;
  assign tile__reset[2] = reset;
  assign tile__clk[3] = clk;
  assign tile__reset[3] = reset;
  assign tile__clk[4] = clk;
  assign tile__reset[4] = reset;
  assign tile__clk[5] = clk;
  assign tile__reset[5] = reset;
  assign tile__clk[6] = clk;
  assign tile__reset[6] = reset;
  assign tile__clk[7] = clk;
  assign tile__reset[7] = reset;
  assign tile__clk[8] = clk;
  assign tile__reset[8] = reset;
  assign tile__clk[9] = clk;
  assign tile__reset[9] = reset;
  assign tile__clk[10] = clk;
  assign tile__reset[10] = reset;
  assign tile__clk[11] = clk;
  assign tile__reset[11] = reset;
  assign tile__clk[12] = clk;
  assign tile__reset[12] = reset;
  assign tile__clk[13] = clk;
  assign tile__reset[13] = reset;
  assign tile__clk[14] = clk;
  assign tile__reset[14] = reset;
  assign tile__clk[15] = clk;
  assign tile__reset[15] = reset;
  assign data_mem__clk = clk;
  assign data_mem__reset = reset;
  assign tile__recv_waddr__en[0] = recv_waddr__en[0];
  assign tile__recv_waddr__msg[0] = recv_waddr__msg[0];
  assign recv_waddr__rdy[0] = tile__recv_waddr__rdy[0];
  assign tile__recv_wopt__en[0] = recv_wopt__en[0];
  assign tile__recv_wopt__msg[0] = recv_wopt__msg[0];
  assign recv_wopt__rdy[0] = tile__recv_wopt__rdy[0];
  assign tile__recv_data__en[4][1] = tile__send_data__en[0][0];
  assign tile__recv_data__msg[4][1] = tile__send_data__msg[0][0];
  assign tile__send_data__rdy[0][0] = tile__recv_data__rdy[4][1];
  assign tile__recv_data__en[1][2] = tile__send_data__en[0][3];
  assign tile__recv_data__msg[1][2] = tile__send_data__msg[0][3];
  assign tile__send_data__rdy[0][3] = tile__recv_data__rdy[1][2];
  assign tile__send_data__rdy[0][1] = 1'd0;
  assign tile__recv_data__en[0][1] = 1'd0;
  assign tile__recv_data__msg[0][1] = { 32'd0, 1'd0, 1'd0 };
  assign tile__send_data__rdy[0][2] = 1'd0;
  assign tile__recv_data__en[0][2] = 1'd0;
  assign tile__recv_data__msg[0][2] = { 32'd0, 1'd0, 1'd0 };
  assign data_mem__recv_raddr__en[0] = tile__to_mem_raddr__en[0];
  assign data_mem__recv_raddr__msg[0] = tile__to_mem_raddr__msg[0];
  assign tile__to_mem_raddr__rdy[0] = data_mem__recv_raddr__rdy[0];
  assign tile__from_mem_rdata__en[0] = data_mem__send_rdata__en[0];
  assign tile__from_mem_rdata__msg[0] = data_mem__send_rdata__msg[0];
  assign data_mem__send_rdata__rdy[0] = tile__from_mem_rdata__rdy[0];
  assign data_mem__recv_waddr__en[0] = tile__to_mem_waddr__en[0];
  assign data_mem__recv_waddr__msg[0] = tile__to_mem_waddr__msg[0];
  assign tile__to_mem_waddr__rdy[0] = data_mem__recv_waddr__rdy[0];
  assign data_mem__recv_wdata__en[0] = tile__to_mem_wdata__en[0];
  assign data_mem__recv_wdata__msg[0] = tile__to_mem_wdata__msg[0];
  assign tile__to_mem_wdata__rdy[0] = data_mem__recv_wdata__rdy[0];
  assign tile__recv_waddr__en[1] = recv_waddr__en[1];
  assign tile__recv_waddr__msg[1] = recv_waddr__msg[1];
  assign recv_waddr__rdy[1] = tile__recv_waddr__rdy[1];
  assign tile__recv_wopt__en[1] = recv_wopt__en[1];
  assign tile__recv_wopt__msg[1] = recv_wopt__msg[1];
  assign recv_wopt__rdy[1] = tile__recv_wopt__rdy[1];
  assign tile__recv_data__en[5][1] = tile__send_data__en[1][0];
  assign tile__recv_data__msg[5][1] = tile__send_data__msg[1][0];
  assign tile__send_data__rdy[1][0] = tile__recv_data__rdy[5][1];
  assign tile__recv_data__en[0][3] = tile__send_data__en[1][2];
  assign tile__recv_data__msg[0][3] = tile__send_data__msg[1][2];
  assign tile__send_data__rdy[1][2] = tile__recv_data__rdy[0][3];
  assign tile__recv_data__en[2][2] = tile__send_data__en[1][3];
  assign tile__recv_data__msg[2][2] = tile__send_data__msg[1][3];
  assign tile__send_data__rdy[1][3] = tile__recv_data__rdy[2][2];
  assign tile__send_data__rdy[1][1] = 1'd0;
  assign tile__recv_data__en[1][1] = 1'd0;
  assign tile__recv_data__msg[1][1] = { 32'd0, 1'd0, 1'd0 };
  assign tile__to_mem_raddr__rdy[1] = 1'd0;
  assign tile__from_mem_rdata__en[1] = 1'd0;
  assign tile__from_mem_rdata__msg[1] = { 32'd0, 1'd0, 1'd0 };
  assign tile__to_mem_waddr__rdy[1] = 1'd0;
  assign tile__to_mem_wdata__rdy[1] = 1'd0;
  assign tile__recv_waddr__en[2] = recv_waddr__en[2];
  assign tile__recv_waddr__msg[2] = recv_waddr__msg[2];
  assign recv_waddr__rdy[2] = tile__recv_waddr__rdy[2];
  assign tile__recv_wopt__en[2] = recv_wopt__en[2];
  assign tile__recv_wopt__msg[2] = recv_wopt__msg[2];
  assign recv_wopt__rdy[2] = tile__recv_wopt__rdy[2];
  assign tile__recv_data__en[6][1] = tile__send_data__en[2][0];
  assign tile__recv_data__msg[6][1] = tile__send_data__msg[2][0];
  assign tile__send_data__rdy[2][0] = tile__recv_data__rdy[6][1];
  assign tile__recv_data__en[1][3] = tile__send_data__en[2][2];
  assign tile__recv_data__msg[1][3] = tile__send_data__msg[2][2];
  assign tile__send_data__rdy[2][2] = tile__recv_data__rdy[1][3];
  assign tile__recv_data__en[3][2] = tile__send_data__en[2][3];
  assign tile__recv_data__msg[3][2] = tile__send_data__msg[2][3];
  assign tile__send_data__rdy[2][3] = tile__recv_data__rdy[3][2];
  assign tile__send_data__rdy[2][1] = 1'd0;
  assign tile__recv_data__en[2][1] = 1'd0;
  assign tile__recv_data__msg[2][1] = { 32'd0, 1'd0, 1'd0 };
  assign tile__to_mem_raddr__rdy[2] = 1'd0;
  assign tile__from_mem_rdata__en[2] = 1'd0;
  assign tile__from_mem_rdata__msg[2] = { 32'd0, 1'd0, 1'd0 };
  assign tile__to_mem_waddr__rdy[2] = 1'd0;
  assign tile__to_mem_wdata__rdy[2] = 1'd0;
  assign tile__recv_waddr__en[3] = recv_waddr__en[3];
  assign tile__recv_waddr__msg[3] = recv_waddr__msg[3];
  assign recv_waddr__rdy[3] = tile__recv_waddr__rdy[3];
  assign tile__recv_wopt__en[3] = recv_wopt__en[3];
  assign tile__recv_wopt__msg[3] = recv_wopt__msg[3];
  assign recv_wopt__rdy[3] = tile__recv_wopt__rdy[3];
  assign tile__recv_data__en[7][1] = tile__send_data__en[3][0];
  assign tile__recv_data__msg[7][1] = tile__send_data__msg[3][0];
  assign tile__send_data__rdy[3][0] = tile__recv_data__rdy[7][1];
  assign tile__recv_data__en[2][3] = tile__send_data__en[3][2];
  assign tile__recv_data__msg[2][3] = tile__send_data__msg[3][2];
  assign tile__send_data__rdy[3][2] = tile__recv_data__rdy[2][3];
  assign tile__send_data__rdy[3][1] = 1'd0;
  assign tile__recv_data__en[3][1] = 1'd0;
  assign tile__recv_data__msg[3][1] = { 32'd0, 1'd0, 1'd0 };
  assign tile__send_data__rdy[3][3] = 1'd0;
  assign tile__recv_data__en[3][3] = 1'd0;
  assign tile__recv_data__msg[3][3] = { 32'd0, 1'd0, 1'd0 };
  assign tile__to_mem_raddr__rdy[3] = 1'd0;
  assign tile__from_mem_rdata__en[3] = 1'd0;
  assign tile__from_mem_rdata__msg[3] = { 32'd0, 1'd0, 1'd0 };
  assign tile__to_mem_waddr__rdy[3] = 1'd0;
  assign tile__to_mem_wdata__rdy[3] = 1'd0;
  assign tile__recv_waddr__en[4] = recv_waddr__en[4];
  assign tile__recv_waddr__msg[4] = recv_waddr__msg[4];
  assign recv_waddr__rdy[4] = tile__recv_waddr__rdy[4];
  assign tile__recv_wopt__en[4] = recv_wopt__en[4];
  assign tile__recv_wopt__msg[4] = recv_wopt__msg[4];
  assign recv_wopt__rdy[4] = tile__recv_wopt__rdy[4];
  assign tile__recv_data__en[0][0] = tile__send_data__en[4][1];
  assign tile__recv_data__msg[0][0] = tile__send_data__msg[4][1];
  assign tile__send_data__rdy[4][1] = tile__recv_data__rdy[0][0];
  assign tile__recv_data__en[8][1] = tile__send_data__en[4][0];
  assign tile__recv_data__msg[8][1] = tile__send_data__msg[4][0];
  assign tile__send_data__rdy[4][0] = tile__recv_data__rdy[8][1];
  assign tile__recv_data__en[5][2] = tile__send_data__en[4][3];
  assign tile__recv_data__msg[5][2] = tile__send_data__msg[4][3];
  assign tile__send_data__rdy[4][3] = tile__recv_data__rdy[5][2];
  assign tile__send_data__rdy[4][2] = 1'd0;
  assign tile__recv_data__en[4][2] = 1'd0;
  assign tile__recv_data__msg[4][2] = { 32'd0, 1'd0, 1'd0 };
  assign data_mem__recv_raddr__en[1] = tile__to_mem_raddr__en[4];
  assign data_mem__recv_raddr__msg[1] = tile__to_mem_raddr__msg[4];
  assign tile__to_mem_raddr__rdy[4] = data_mem__recv_raddr__rdy[1];
  assign tile__from_mem_rdata__en[4] = data_mem__send_rdata__en[1];
  assign tile__from_mem_rdata__msg[4] = data_mem__send_rdata__msg[1];
  assign data_mem__send_rdata__rdy[1] = tile__from_mem_rdata__rdy[4];
  assign data_mem__recv_waddr__en[1] = tile__to_mem_waddr__en[4];
  assign data_mem__recv_waddr__msg[1] = tile__to_mem_waddr__msg[4];
  assign tile__to_mem_waddr__rdy[4] = data_mem__recv_waddr__rdy[1];
  assign data_mem__recv_wdata__en[1] = tile__to_mem_wdata__en[4];
  assign data_mem__recv_wdata__msg[1] = tile__to_mem_wdata__msg[4];
  assign tile__to_mem_wdata__rdy[4] = data_mem__recv_wdata__rdy[1];
  assign tile__recv_waddr__en[5] = recv_waddr__en[5];
  assign tile__recv_waddr__msg[5] = recv_waddr__msg[5];
  assign recv_waddr__rdy[5] = tile__recv_waddr__rdy[5];
  assign tile__recv_wopt__en[5] = recv_wopt__en[5];
  assign tile__recv_wopt__msg[5] = recv_wopt__msg[5];
  assign recv_wopt__rdy[5] = tile__recv_wopt__rdy[5];
  assign tile__recv_data__en[1][0] = tile__send_data__en[5][1];
  assign tile__recv_data__msg[1][0] = tile__send_data__msg[5][1];
  assign tile__send_data__rdy[5][1] = tile__recv_data__rdy[1][0];
  assign tile__recv_data__en[9][1] = tile__send_data__en[5][0];
  assign tile__recv_data__msg[9][1] = tile__send_data__msg[5][0];
  assign tile__send_data__rdy[5][0] = tile__recv_data__rdy[9][1];
  assign tile__recv_data__en[4][3] = tile__send_data__en[5][2];
  assign tile__recv_data__msg[4][3] = tile__send_data__msg[5][2];
  assign tile__send_data__rdy[5][2] = tile__recv_data__rdy[4][3];
  assign tile__recv_data__en[6][2] = tile__send_data__en[5][3];
  assign tile__recv_data__msg[6][2] = tile__send_data__msg[5][3];
  assign tile__send_data__rdy[5][3] = tile__recv_data__rdy[6][2];
  assign tile__to_mem_raddr__rdy[5] = 1'd0;
  assign tile__from_mem_rdata__en[5] = 1'd0;
  assign tile__from_mem_rdata__msg[5] = { 32'd0, 1'd0, 1'd0 };
  assign tile__to_mem_waddr__rdy[5] = 1'd0;
  assign tile__to_mem_wdata__rdy[5] = 1'd0;
  assign tile__recv_waddr__en[6] = recv_waddr__en[6];
  assign tile__recv_waddr__msg[6] = recv_waddr__msg[6];
  assign recv_waddr__rdy[6] = tile__recv_waddr__rdy[6];
  assign tile__recv_wopt__en[6] = recv_wopt__en[6];
  assign tile__recv_wopt__msg[6] = recv_wopt__msg[6];
  assign recv_wopt__rdy[6] = tile__recv_wopt__rdy[6];
  assign tile__recv_data__en[2][0] = tile__send_data__en[6][1];
  assign tile__recv_data__msg[2][0] = tile__send_data__msg[6][1];
  assign tile__send_data__rdy[6][1] = tile__recv_data__rdy[2][0];
  assign tile__recv_data__en[10][1] = tile__send_data__en[6][0];
  assign tile__recv_data__msg[10][1] = tile__send_data__msg[6][0];
  assign tile__send_data__rdy[6][0] = tile__recv_data__rdy[10][1];
  assign tile__recv_data__en[5][3] = tile__send_data__en[6][2];
  assign tile__recv_data__msg[5][3] = tile__send_data__msg[6][2];
  assign tile__send_data__rdy[6][2] = tile__recv_data__rdy[5][3];
  assign tile__recv_data__en[7][2] = tile__send_data__en[6][3];
  assign tile__recv_data__msg[7][2] = tile__send_data__msg[6][3];
  assign tile__send_data__rdy[6][3] = tile__recv_data__rdy[7][2];
  assign tile__to_mem_raddr__rdy[6] = 1'd0;
  assign tile__from_mem_rdata__en[6] = 1'd0;
  assign tile__from_mem_rdata__msg[6] = { 32'd0, 1'd0, 1'd0 };
  assign tile__to_mem_waddr__rdy[6] = 1'd0;
  assign tile__to_mem_wdata__rdy[6] = 1'd0;
  assign tile__recv_waddr__en[7] = recv_waddr__en[7];
  assign tile__recv_waddr__msg[7] = recv_waddr__msg[7];
  assign recv_waddr__rdy[7] = tile__recv_waddr__rdy[7];
  assign tile__recv_wopt__en[7] = recv_wopt__en[7];
  assign tile__recv_wopt__msg[7] = recv_wopt__msg[7];
  assign recv_wopt__rdy[7] = tile__recv_wopt__rdy[7];
  assign tile__recv_data__en[3][0] = tile__send_data__en[7][1];
  assign tile__recv_data__msg[3][0] = tile__send_data__msg[7][1];
  assign tile__send_data__rdy[7][1] = tile__recv_data__rdy[3][0];
  assign tile__recv_data__en[11][1] = tile__send_data__en[7][0];
  assign tile__recv_data__msg[11][1] = tile__send_data__msg[7][0];
  assign tile__send_data__rdy[7][0] = tile__recv_data__rdy[11][1];
  assign tile__recv_data__en[6][3] = tile__send_data__en[7][2];
  assign tile__recv_data__msg[6][3] = tile__send_data__msg[7][2];
  assign tile__send_data__rdy[7][2] = tile__recv_data__rdy[6][3];
  assign tile__send_data__rdy[7][3] = 1'd0;
  assign tile__recv_data__en[7][3] = 1'd0;
  assign tile__recv_data__msg[7][3] = { 32'd0, 1'd0, 1'd0 };
  assign tile__to_mem_raddr__rdy[7] = 1'd0;
  assign tile__from_mem_rdata__en[7] = 1'd0;
  assign tile__from_mem_rdata__msg[7] = { 32'd0, 1'd0, 1'd0 };
  assign tile__to_mem_waddr__rdy[7] = 1'd0;
  assign tile__to_mem_wdata__rdy[7] = 1'd0;
  assign tile__recv_waddr__en[8] = recv_waddr__en[8];
  assign tile__recv_waddr__msg[8] = recv_waddr__msg[8];
  assign recv_waddr__rdy[8] = tile__recv_waddr__rdy[8];
  assign tile__recv_wopt__en[8] = recv_wopt__en[8];
  assign tile__recv_wopt__msg[8] = recv_wopt__msg[8];
  assign recv_wopt__rdy[8] = tile__recv_wopt__rdy[8];
  assign tile__recv_data__en[4][0] = tile__send_data__en[8][1];
  assign tile__recv_data__msg[4][0] = tile__send_data__msg[8][1];
  assign tile__send_data__rdy[8][1] = tile__recv_data__rdy[4][0];
  assign tile__recv_data__en[12][1] = tile__send_data__en[8][0];
  assign tile__recv_data__msg[12][1] = tile__send_data__msg[8][0];
  assign tile__send_data__rdy[8][0] = tile__recv_data__rdy[12][1];
  assign tile__recv_data__en[9][2] = tile__send_data__en[8][3];
  assign tile__recv_data__msg[9][2] = tile__send_data__msg[8][3];
  assign tile__send_data__rdy[8][3] = tile__recv_data__rdy[9][2];
  assign tile__send_data__rdy[8][2] = 1'd0;
  assign tile__recv_data__en[8][2] = 1'd0;
  assign tile__recv_data__msg[8][2] = { 32'd0, 1'd0, 1'd0 };
  assign data_mem__recv_raddr__en[2] = tile__to_mem_raddr__en[8];
  assign data_mem__recv_raddr__msg[2] = tile__to_mem_raddr__msg[8];
  assign tile__to_mem_raddr__rdy[8] = data_mem__recv_raddr__rdy[2];
  assign tile__from_mem_rdata__en[8] = data_mem__send_rdata__en[2];
  assign tile__from_mem_rdata__msg[8] = data_mem__send_rdata__msg[2];
  assign data_mem__send_rdata__rdy[2] = tile__from_mem_rdata__rdy[8];
  assign data_mem__recv_waddr__en[2] = tile__to_mem_waddr__en[8];
  assign data_mem__recv_waddr__msg[2] = tile__to_mem_waddr__msg[8];
  assign tile__to_mem_waddr__rdy[8] = data_mem__recv_waddr__rdy[2];
  assign data_mem__recv_wdata__en[2] = tile__to_mem_wdata__en[8];
  assign data_mem__recv_wdata__msg[2] = tile__to_mem_wdata__msg[8];
  assign tile__to_mem_wdata__rdy[8] = data_mem__recv_wdata__rdy[2];
  assign tile__recv_waddr__en[9] = recv_waddr__en[9];
  assign tile__recv_waddr__msg[9] = recv_waddr__msg[9];
  assign recv_waddr__rdy[9] = tile__recv_waddr__rdy[9];
  assign tile__recv_wopt__en[9] = recv_wopt__en[9];
  assign tile__recv_wopt__msg[9] = recv_wopt__msg[9];
  assign recv_wopt__rdy[9] = tile__recv_wopt__rdy[9];
  assign tile__recv_data__en[5][0] = tile__send_data__en[9][1];
  assign tile__recv_data__msg[5][0] = tile__send_data__msg[9][1];
  assign tile__send_data__rdy[9][1] = tile__recv_data__rdy[5][0];
  assign tile__recv_data__en[13][1] = tile__send_data__en[9][0];
  assign tile__recv_data__msg[13][1] = tile__send_data__msg[9][0];
  assign tile__send_data__rdy[9][0] = tile__recv_data__rdy[13][1];
  assign tile__recv_data__en[8][3] = tile__send_data__en[9][2];
  assign tile__recv_data__msg[8][3] = tile__send_data__msg[9][2];
  assign tile__send_data__rdy[9][2] = tile__recv_data__rdy[8][3];
  assign tile__recv_data__en[10][2] = tile__send_data__en[9][3];
  assign tile__recv_data__msg[10][2] = tile__send_data__msg[9][3];
  assign tile__send_data__rdy[9][3] = tile__recv_data__rdy[10][2];
  assign tile__to_mem_raddr__rdy[9] = 1'd0;
  assign tile__from_mem_rdata__en[9] = 1'd0;
  assign tile__from_mem_rdata__msg[9] = { 32'd0, 1'd0, 1'd0 };
  assign tile__to_mem_waddr__rdy[9] = 1'd0;
  assign tile__to_mem_wdata__rdy[9] = 1'd0;
  assign tile__recv_waddr__en[10] = recv_waddr__en[10];
  assign tile__recv_waddr__msg[10] = recv_waddr__msg[10];
  assign recv_waddr__rdy[10] = tile__recv_waddr__rdy[10];
  assign tile__recv_wopt__en[10] = recv_wopt__en[10];
  assign tile__recv_wopt__msg[10] = recv_wopt__msg[10];
  assign recv_wopt__rdy[10] = tile__recv_wopt__rdy[10];
  assign tile__recv_data__en[6][0] = tile__send_data__en[10][1];
  assign tile__recv_data__msg[6][0] = tile__send_data__msg[10][1];
  assign tile__send_data__rdy[10][1] = tile__recv_data__rdy[6][0];
  assign tile__recv_data__en[14][1] = tile__send_data__en[10][0];
  assign tile__recv_data__msg[14][1] = tile__send_data__msg[10][0];
  assign tile__send_data__rdy[10][0] = tile__recv_data__rdy[14][1];
  assign tile__recv_data__en[9][3] = tile__send_data__en[10][2];
  assign tile__recv_data__msg[9][3] = tile__send_data__msg[10][2];
  assign tile__send_data__rdy[10][2] = tile__recv_data__rdy[9][3];
  assign tile__recv_data__en[11][2] = tile__send_data__en[10][3];
  assign tile__recv_data__msg[11][2] = tile__send_data__msg[10][3];
  assign tile__send_data__rdy[10][3] = tile__recv_data__rdy[11][2];
  assign tile__to_mem_raddr__rdy[10] = 1'd0;
  assign tile__from_mem_rdata__en[10] = 1'd0;
  assign tile__from_mem_rdata__msg[10] = { 32'd0, 1'd0, 1'd0 };
  assign tile__to_mem_waddr__rdy[10] = 1'd0;
  assign tile__to_mem_wdata__rdy[10] = 1'd0;
  assign tile__recv_waddr__en[11] = recv_waddr__en[11];
  assign tile__recv_waddr__msg[11] = recv_waddr__msg[11];
  assign recv_waddr__rdy[11] = tile__recv_waddr__rdy[11];
  assign tile__recv_wopt__en[11] = recv_wopt__en[11];
  assign tile__recv_wopt__msg[11] = recv_wopt__msg[11];
  assign recv_wopt__rdy[11] = tile__recv_wopt__rdy[11];
  assign tile__recv_data__en[7][0] = tile__send_data__en[11][1];
  assign tile__recv_data__msg[7][0] = tile__send_data__msg[11][1];
  assign tile__send_data__rdy[11][1] = tile__recv_data__rdy[7][0];
  assign tile__recv_data__en[15][1] = tile__send_data__en[11][0];
  assign tile__recv_data__msg[15][1] = tile__send_data__msg[11][0];
  assign tile__send_data__rdy[11][0] = tile__recv_data__rdy[15][1];
  assign tile__recv_data__en[10][3] = tile__send_data__en[11][2];
  assign tile__recv_data__msg[10][3] = tile__send_data__msg[11][2];
  assign tile__send_data__rdy[11][2] = tile__recv_data__rdy[10][3];
  assign tile__send_data__rdy[11][3] = 1'd0;
  assign tile__recv_data__en[11][3] = 1'd0;
  assign tile__recv_data__msg[11][3] = { 32'd0, 1'd0, 1'd0 };
  assign tile__to_mem_raddr__rdy[11] = 1'd0;
  assign tile__from_mem_rdata__en[11] = 1'd0;
  assign tile__from_mem_rdata__msg[11] = { 32'd0, 1'd0, 1'd0 };
  assign tile__to_mem_waddr__rdy[11] = 1'd0;
  assign tile__to_mem_wdata__rdy[11] = 1'd0;
  assign tile__recv_waddr__en[12] = recv_waddr__en[12];
  assign tile__recv_waddr__msg[12] = recv_waddr__msg[12];
  assign recv_waddr__rdy[12] = tile__recv_waddr__rdy[12];
  assign tile__recv_wopt__en[12] = recv_wopt__en[12];
  assign tile__recv_wopt__msg[12] = recv_wopt__msg[12];
  assign recv_wopt__rdy[12] = tile__recv_wopt__rdy[12];
  assign tile__recv_data__en[8][0] = tile__send_data__en[12][1];
  assign tile__recv_data__msg[8][0] = tile__send_data__msg[12][1];
  assign tile__send_data__rdy[12][1] = tile__recv_data__rdy[8][0];
  assign tile__recv_data__en[13][2] = tile__send_data__en[12][3];
  assign tile__recv_data__msg[13][2] = tile__send_data__msg[12][3];
  assign tile__send_data__rdy[12][3] = tile__recv_data__rdy[13][2];
  assign tile__send_data__rdy[12][0] = 1'd0;
  assign tile__recv_data__en[12][0] = 1'd0;
  assign tile__recv_data__msg[12][0] = { 32'd0, 1'd0, 1'd0 };
  assign tile__send_data__rdy[12][2] = 1'd0;
  assign tile__recv_data__en[12][2] = 1'd0;
  assign tile__recv_data__msg[12][2] = { 32'd0, 1'd0, 1'd0 };
  assign data_mem__recv_raddr__en[3] = tile__to_mem_raddr__en[12];
  assign data_mem__recv_raddr__msg[3] = tile__to_mem_raddr__msg[12];
  assign tile__to_mem_raddr__rdy[12] = data_mem__recv_raddr__rdy[3];
  assign tile__from_mem_rdata__en[12] = data_mem__send_rdata__en[3];
  assign tile__from_mem_rdata__msg[12] = data_mem__send_rdata__msg[3];
  assign data_mem__send_rdata__rdy[3] = tile__from_mem_rdata__rdy[12];
  assign data_mem__recv_waddr__en[3] = tile__to_mem_waddr__en[12];
  assign data_mem__recv_waddr__msg[3] = tile__to_mem_waddr__msg[12];
  assign tile__to_mem_waddr__rdy[12] = data_mem__recv_waddr__rdy[3];
  assign data_mem__recv_wdata__en[3] = tile__to_mem_wdata__en[12];
  assign data_mem__recv_wdata__msg[3] = tile__to_mem_wdata__msg[12];
  assign tile__to_mem_wdata__rdy[12] = data_mem__recv_wdata__rdy[3];
  assign tile__recv_waddr__en[13] = recv_waddr__en[13];
  assign tile__recv_waddr__msg[13] = recv_waddr__msg[13];
  assign recv_waddr__rdy[13] = tile__recv_waddr__rdy[13];
  assign tile__recv_wopt__en[13] = recv_wopt__en[13];
  assign tile__recv_wopt__msg[13] = recv_wopt__msg[13];
  assign recv_wopt__rdy[13] = tile__recv_wopt__rdy[13];
  assign tile__recv_data__en[9][0] = tile__send_data__en[13][1];
  assign tile__recv_data__msg[9][0] = tile__send_data__msg[13][1];
  assign tile__send_data__rdy[13][1] = tile__recv_data__rdy[9][0];
  assign tile__recv_data__en[12][3] = tile__send_data__en[13][2];
  assign tile__recv_data__msg[12][3] = tile__send_data__msg[13][2];
  assign tile__send_data__rdy[13][2] = tile__recv_data__rdy[12][3];
  assign tile__recv_data__en[14][2] = tile__send_data__en[13][3];
  assign tile__recv_data__msg[14][2] = tile__send_data__msg[13][3];
  assign tile__send_data__rdy[13][3] = tile__recv_data__rdy[14][2];
  assign tile__send_data__rdy[13][0] = 1'd0;
  assign tile__recv_data__en[13][0] = 1'd0;
  assign tile__recv_data__msg[13][0] = { 32'd0, 1'd0, 1'd0 };
  assign tile__to_mem_raddr__rdy[13] = 1'd0;
  assign tile__from_mem_rdata__en[13] = 1'd0;
  assign tile__from_mem_rdata__msg[13] = { 32'd0, 1'd0, 1'd0 };
  assign tile__to_mem_waddr__rdy[13] = 1'd0;
  assign tile__to_mem_wdata__rdy[13] = 1'd0;
  assign tile__recv_waddr__en[14] = recv_waddr__en[14];
  assign tile__recv_waddr__msg[14] = recv_waddr__msg[14];
  assign recv_waddr__rdy[14] = tile__recv_waddr__rdy[14];
  assign tile__recv_wopt__en[14] = recv_wopt__en[14];
  assign tile__recv_wopt__msg[14] = recv_wopt__msg[14];
  assign recv_wopt__rdy[14] = tile__recv_wopt__rdy[14];
  assign tile__recv_data__en[10][0] = tile__send_data__en[14][1];
  assign tile__recv_data__msg[10][0] = tile__send_data__msg[14][1];
  assign tile__send_data__rdy[14][1] = tile__recv_data__rdy[10][0];
  assign tile__recv_data__en[13][3] = tile__send_data__en[14][2];
  assign tile__recv_data__msg[13][3] = tile__send_data__msg[14][2];
  assign tile__send_data__rdy[14][2] = tile__recv_data__rdy[13][3];
  assign tile__recv_data__en[15][2] = tile__send_data__en[14][3];
  assign tile__recv_data__msg[15][2] = tile__send_data__msg[14][3];
  assign tile__send_data__rdy[14][3] = tile__recv_data__rdy[15][2];
  assign tile__send_data__rdy[14][0] = 1'd0;
  assign tile__recv_data__en[14][0] = 1'd0;
  assign tile__recv_data__msg[14][0] = { 32'd0, 1'd0, 1'd0 };
  assign tile__to_mem_raddr__rdy[14] = 1'd0;
  assign tile__from_mem_rdata__en[14] = 1'd0;
  assign tile__from_mem_rdata__msg[14] = { 32'd0, 1'd0, 1'd0 };
  assign tile__to_mem_waddr__rdy[14] = 1'd0;
  assign tile__to_mem_wdata__rdy[14] = 1'd0;
  assign tile__recv_waddr__en[15] = recv_waddr__en[15];
  assign tile__recv_waddr__msg[15] = recv_waddr__msg[15];
  assign recv_waddr__rdy[15] = tile__recv_waddr__rdy[15];
  assign tile__recv_wopt__en[15] = recv_wopt__en[15];
  assign tile__recv_wopt__msg[15] = recv_wopt__msg[15];
  assign recv_wopt__rdy[15] = tile__recv_wopt__rdy[15];
  assign tile__recv_data__en[11][0] = tile__send_data__en[15][1];
  assign tile__recv_data__msg[11][0] = tile__send_data__msg[15][1];
  assign tile__send_data__rdy[15][1] = tile__recv_data__rdy[11][0];
  assign tile__recv_data__en[14][3] = tile__send_data__en[15][2];
  assign tile__recv_data__msg[14][3] = tile__send_data__msg[15][2];
  assign tile__send_data__rdy[15][2] = tile__recv_data__rdy[14][3];
  assign tile__send_data__rdy[15][0] = 1'd0;
  assign tile__recv_data__en[15][0] = 1'd0;
  assign tile__recv_data__msg[15][0] = { 32'd0, 1'd0, 1'd0 };
  assign tile__send_data__rdy[15][3] = 1'd0;
  assign tile__recv_data__en[15][3] = 1'd0;
  assign tile__recv_data__msg[15][3] = { 32'd0, 1'd0, 1'd0 };
  assign tile__to_mem_raddr__rdy[15] = 1'd0;
  assign tile__from_mem_rdata__en[15] = 1'd0;
  assign tile__from_mem_rdata__msg[15] = { 32'd0, 1'd0, 1'd0 };
  assign tile__to_mem_waddr__rdy[15] = 1'd0;
  assign tile__to_mem_wdata__rdy[15] = 1'd0;

endmodule
